library verilog;
use verilog.vl_types.all;
entity Acumulador_vlg_check_tst is
    port(
        AC_out          : in     vl_logic_vector(15 downto 0);
        sampler_rx      : in     vl_logic
    );
end Acumulador_vlg_check_tst;
