library verilog;
use verilog.vl_types.all;
entity OperatorMUX_vlg_vec_tst is
end OperatorMUX_vlg_vec_tst;
