library verilog;
use verilog.vl_types.all;
entity Data_MdMux_vlg_vec_tst is
end Data_MdMux_vlg_vec_tst;
