library verilog;
use verilog.vl_types.all;
entity GeneralPR_vlg_vec_tst is
end GeneralPR_vlg_vec_tst;
