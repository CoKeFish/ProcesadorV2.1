library verilog;
use verilog.vl_types.all;
entity DirMdMux_vlg_vec_tst is
end DirMdMux_vlg_vec_tst;
