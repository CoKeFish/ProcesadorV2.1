library verilog;
use verilog.vl_types.all;
entity ProgramCounterMUX_vlg_vec_tst is
end ProgramCounterMUX_vlg_vec_tst;
