library verilog;
use verilog.vl_types.all;
entity AcumMUX_vlg_vec_tst is
end AcumMUX_vlg_vec_tst;
