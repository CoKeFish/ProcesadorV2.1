library verilog;
use verilog.vl_types.all;
entity Computador_vlg_vec_tst is
end Computador_vlg_vec_tst;
