library verilog;
use verilog.vl_types.all;
entity DirRegister_vlg_vec_tst is
end DirRegister_vlg_vec_tst;
