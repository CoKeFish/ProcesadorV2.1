library verilog;
use verilog.vl_types.all;
entity ProgramStatus_vlg_vec_tst is
end ProgramStatus_vlg_vec_tst;
