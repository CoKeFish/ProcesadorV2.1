library verilog;
use verilog.vl_types.all;
entity StackPointer_vlg_vec_tst is
end StackPointer_vlg_vec_tst;
