library verilog;
use verilog.vl_types.all;
entity Acumulador_vlg_vec_tst is
end Acumulador_vlg_vec_tst;
