library verilog;
use verilog.vl_types.all;
entity AcumMux_vlg_vec_tst is
end AcumMux_vlg_vec_tst;
