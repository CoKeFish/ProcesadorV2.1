library verilog;
use verilog.vl_types.all;
entity PSRMux_vlg_vec_tst is
end PSRMux_vlg_vec_tst;
