library verilog;
use verilog.vl_types.all;
entity ALUMux_vlg_vec_tst is
end ALUMux_vlg_vec_tst;
